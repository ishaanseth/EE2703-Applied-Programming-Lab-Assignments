.circuit
V1 N1 0 DC 5
R1 N1 N2 1k
.end
